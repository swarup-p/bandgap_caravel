magic
tech sky130A
timestamp 1616700505
<< mvnmos >>
rect 225 601 825 4801
<< mvndiff >>
rect 190 4768 225 4801
rect 190 4750 199 4768
rect 216 4750 225 4768
rect 190 4732 225 4750
rect 190 4714 199 4732
rect 216 4714 225 4732
rect 190 4696 225 4714
rect 190 4678 199 4696
rect 216 4678 225 4696
rect 190 4660 225 4678
rect 190 4642 199 4660
rect 216 4642 225 4660
rect 190 4624 225 4642
rect 190 4606 199 4624
rect 216 4606 225 4624
rect 190 4588 225 4606
rect 190 4570 199 4588
rect 216 4570 225 4588
rect 190 4552 225 4570
rect 190 4534 199 4552
rect 216 4534 225 4552
rect 190 4516 225 4534
rect 190 4498 199 4516
rect 216 4498 225 4516
rect 190 4480 225 4498
rect 190 4462 199 4480
rect 216 4462 225 4480
rect 190 4444 225 4462
rect 190 4426 199 4444
rect 216 4426 225 4444
rect 190 4408 225 4426
rect 190 4390 199 4408
rect 216 4390 225 4408
rect 190 4372 225 4390
rect 190 4354 199 4372
rect 216 4354 225 4372
rect 190 4336 225 4354
rect 190 4318 199 4336
rect 216 4318 225 4336
rect 190 4300 225 4318
rect 190 4282 199 4300
rect 216 4282 225 4300
rect 190 4264 225 4282
rect 190 4246 199 4264
rect 216 4246 225 4264
rect 190 4228 225 4246
rect 190 4210 199 4228
rect 216 4210 225 4228
rect 190 4192 225 4210
rect 190 4174 199 4192
rect 216 4174 225 4192
rect 190 4156 225 4174
rect 190 4138 199 4156
rect 216 4138 225 4156
rect 190 4120 225 4138
rect 190 4102 199 4120
rect 216 4102 225 4120
rect 190 4084 225 4102
rect 190 4066 199 4084
rect 216 4066 225 4084
rect 190 4048 225 4066
rect 190 4030 199 4048
rect 216 4030 225 4048
rect 190 4012 225 4030
rect 190 3994 199 4012
rect 216 3994 225 4012
rect 190 3976 225 3994
rect 190 3958 199 3976
rect 216 3958 225 3976
rect 190 3940 225 3958
rect 190 3922 199 3940
rect 216 3922 225 3940
rect 190 3904 225 3922
rect 190 3886 199 3904
rect 216 3886 225 3904
rect 190 3868 225 3886
rect 190 3850 199 3868
rect 216 3850 225 3868
rect 190 3832 225 3850
rect 190 3814 199 3832
rect 216 3814 225 3832
rect 190 3796 225 3814
rect 190 3778 199 3796
rect 216 3778 225 3796
rect 190 3760 225 3778
rect 190 3742 199 3760
rect 216 3742 225 3760
rect 190 3724 225 3742
rect 190 3706 199 3724
rect 216 3706 225 3724
rect 190 3688 225 3706
rect 190 3670 199 3688
rect 216 3670 225 3688
rect 190 3652 225 3670
rect 190 3634 199 3652
rect 216 3634 225 3652
rect 190 3616 225 3634
rect 190 3598 199 3616
rect 216 3598 225 3616
rect 190 3580 225 3598
rect 190 3562 199 3580
rect 216 3562 225 3580
rect 190 3544 225 3562
rect 190 3526 199 3544
rect 216 3526 225 3544
rect 190 3508 225 3526
rect 190 3490 199 3508
rect 216 3490 225 3508
rect 190 3472 225 3490
rect 190 3454 199 3472
rect 216 3454 225 3472
rect 190 3436 225 3454
rect 190 3418 199 3436
rect 216 3418 225 3436
rect 190 3400 225 3418
rect 190 3382 199 3400
rect 216 3382 225 3400
rect 190 3364 225 3382
rect 190 3346 199 3364
rect 216 3346 225 3364
rect 190 3328 225 3346
rect 190 3310 199 3328
rect 216 3310 225 3328
rect 190 3292 225 3310
rect 190 3274 199 3292
rect 216 3274 225 3292
rect 190 3256 225 3274
rect 190 3238 199 3256
rect 216 3238 225 3256
rect 190 3220 225 3238
rect 190 3202 199 3220
rect 216 3202 225 3220
rect 190 3184 225 3202
rect 190 3166 199 3184
rect 216 3166 225 3184
rect 190 3148 225 3166
rect 190 3130 199 3148
rect 216 3130 225 3148
rect 190 3112 225 3130
rect 190 3094 199 3112
rect 216 3094 225 3112
rect 190 3076 225 3094
rect 190 3058 199 3076
rect 216 3058 225 3076
rect 190 3040 225 3058
rect 190 3022 199 3040
rect 216 3022 225 3040
rect 190 3004 225 3022
rect 190 2986 199 3004
rect 216 2986 225 3004
rect 190 2968 225 2986
rect 190 2950 199 2968
rect 216 2950 225 2968
rect 190 2932 225 2950
rect 190 2914 199 2932
rect 216 2914 225 2932
rect 190 2896 225 2914
rect 190 2878 199 2896
rect 216 2878 225 2896
rect 190 2860 225 2878
rect 190 2842 199 2860
rect 216 2842 225 2860
rect 190 2824 225 2842
rect 190 2806 199 2824
rect 216 2806 225 2824
rect 190 2788 225 2806
rect 190 2770 199 2788
rect 216 2770 225 2788
rect 190 2752 225 2770
rect 190 2734 199 2752
rect 216 2734 225 2752
rect 190 2716 225 2734
rect 190 2698 199 2716
rect 216 2698 225 2716
rect 190 2680 225 2698
rect 190 2662 199 2680
rect 216 2662 225 2680
rect 190 2644 225 2662
rect 190 2626 199 2644
rect 216 2626 225 2644
rect 190 2608 225 2626
rect 190 2590 199 2608
rect 216 2590 225 2608
rect 190 2572 225 2590
rect 190 2554 199 2572
rect 216 2554 225 2572
rect 190 2536 225 2554
rect 190 2518 199 2536
rect 216 2518 225 2536
rect 190 2500 225 2518
rect 190 2482 199 2500
rect 216 2482 225 2500
rect 190 2464 225 2482
rect 190 2446 199 2464
rect 216 2446 225 2464
rect 190 2428 225 2446
rect 190 2410 199 2428
rect 216 2410 225 2428
rect 190 2392 225 2410
rect 190 2374 199 2392
rect 216 2374 225 2392
rect 190 2356 225 2374
rect 190 2338 199 2356
rect 216 2338 225 2356
rect 190 2320 225 2338
rect 190 2302 199 2320
rect 216 2302 225 2320
rect 190 2284 225 2302
rect 190 2266 199 2284
rect 216 2266 225 2284
rect 190 2248 225 2266
rect 190 2230 199 2248
rect 216 2230 225 2248
rect 190 2212 225 2230
rect 190 2194 199 2212
rect 216 2194 225 2212
rect 190 2176 225 2194
rect 190 2158 199 2176
rect 216 2158 225 2176
rect 190 2140 225 2158
rect 190 2122 199 2140
rect 216 2122 225 2140
rect 190 2104 225 2122
rect 190 2086 199 2104
rect 216 2086 225 2104
rect 190 2068 225 2086
rect 190 2050 199 2068
rect 216 2050 225 2068
rect 190 2032 225 2050
rect 190 2014 199 2032
rect 216 2014 225 2032
rect 190 1996 225 2014
rect 190 1978 199 1996
rect 216 1978 225 1996
rect 190 1960 225 1978
rect 190 1942 199 1960
rect 216 1942 225 1960
rect 190 1924 225 1942
rect 190 1906 199 1924
rect 216 1906 225 1924
rect 190 1888 225 1906
rect 190 1870 199 1888
rect 216 1870 225 1888
rect 190 1852 225 1870
rect 190 1834 199 1852
rect 216 1834 225 1852
rect 190 1816 225 1834
rect 190 1798 199 1816
rect 216 1798 225 1816
rect 190 1780 225 1798
rect 190 1762 199 1780
rect 216 1762 225 1780
rect 190 1744 225 1762
rect 190 1726 199 1744
rect 216 1726 225 1744
rect 190 1708 225 1726
rect 190 1690 199 1708
rect 216 1690 225 1708
rect 190 1672 225 1690
rect 190 1654 199 1672
rect 216 1654 225 1672
rect 190 1636 225 1654
rect 190 1618 199 1636
rect 216 1618 225 1636
rect 190 1600 225 1618
rect 190 1582 199 1600
rect 216 1582 225 1600
rect 190 1564 225 1582
rect 190 1546 199 1564
rect 216 1546 225 1564
rect 190 1528 225 1546
rect 190 1510 199 1528
rect 216 1510 225 1528
rect 190 1492 225 1510
rect 190 1474 199 1492
rect 216 1474 225 1492
rect 190 1456 225 1474
rect 190 1438 199 1456
rect 216 1438 225 1456
rect 190 1420 225 1438
rect 190 1402 199 1420
rect 216 1402 225 1420
rect 190 1384 225 1402
rect 190 1366 199 1384
rect 216 1366 225 1384
rect 190 1348 225 1366
rect 190 1330 199 1348
rect 216 1330 225 1348
rect 190 1312 225 1330
rect 190 1294 199 1312
rect 216 1294 225 1312
rect 190 1276 225 1294
rect 190 1258 199 1276
rect 216 1258 225 1276
rect 190 1240 225 1258
rect 190 1222 199 1240
rect 216 1222 225 1240
rect 190 1204 225 1222
rect 190 1186 199 1204
rect 216 1186 225 1204
rect 190 1168 225 1186
rect 190 1150 199 1168
rect 216 1150 225 1168
rect 190 1132 225 1150
rect 190 1114 199 1132
rect 216 1114 225 1132
rect 190 1096 225 1114
rect 190 1078 199 1096
rect 216 1078 225 1096
rect 190 1060 225 1078
rect 190 1042 199 1060
rect 216 1042 225 1060
rect 190 1024 225 1042
rect 190 1006 199 1024
rect 216 1006 225 1024
rect 190 988 225 1006
rect 190 970 199 988
rect 216 970 225 988
rect 190 952 225 970
rect 190 934 199 952
rect 216 934 225 952
rect 190 916 225 934
rect 190 898 199 916
rect 216 898 225 916
rect 190 880 225 898
rect 190 862 199 880
rect 216 862 225 880
rect 190 844 225 862
rect 190 826 199 844
rect 216 826 225 844
rect 190 808 225 826
rect 190 790 199 808
rect 216 790 225 808
rect 190 772 225 790
rect 190 754 199 772
rect 216 754 225 772
rect 190 736 225 754
rect 190 718 199 736
rect 216 718 225 736
rect 190 700 225 718
rect 190 682 199 700
rect 216 682 225 700
rect 190 664 225 682
rect 190 646 199 664
rect 216 646 225 664
rect 190 628 225 646
rect 190 610 199 628
rect 216 610 225 628
rect 190 601 225 610
rect 825 4768 860 4801
rect 825 4750 834 4768
rect 851 4750 860 4768
rect 825 4732 860 4750
rect 825 4714 834 4732
rect 851 4714 860 4732
rect 825 4696 860 4714
rect 825 4678 834 4696
rect 851 4678 860 4696
rect 825 4660 860 4678
rect 825 4642 834 4660
rect 851 4642 860 4660
rect 825 4624 860 4642
rect 825 4606 834 4624
rect 851 4606 860 4624
rect 825 4588 860 4606
rect 825 4570 834 4588
rect 851 4570 860 4588
rect 825 4552 860 4570
rect 825 4534 834 4552
rect 851 4534 860 4552
rect 825 4516 860 4534
rect 825 4498 834 4516
rect 851 4498 860 4516
rect 825 4480 860 4498
rect 825 4462 834 4480
rect 851 4462 860 4480
rect 825 4444 860 4462
rect 825 4426 834 4444
rect 851 4426 860 4444
rect 825 4408 860 4426
rect 825 4390 834 4408
rect 851 4390 860 4408
rect 825 4372 860 4390
rect 825 4354 834 4372
rect 851 4354 860 4372
rect 825 4336 860 4354
rect 825 4318 834 4336
rect 851 4318 860 4336
rect 825 4300 860 4318
rect 825 4282 834 4300
rect 851 4282 860 4300
rect 825 4264 860 4282
rect 825 4246 834 4264
rect 851 4246 860 4264
rect 825 4228 860 4246
rect 825 4210 834 4228
rect 851 4210 860 4228
rect 825 4192 860 4210
rect 825 4174 834 4192
rect 851 4174 860 4192
rect 825 4156 860 4174
rect 825 4138 834 4156
rect 851 4138 860 4156
rect 825 4120 860 4138
rect 825 4102 834 4120
rect 851 4102 860 4120
rect 825 4084 860 4102
rect 825 4066 834 4084
rect 851 4066 860 4084
rect 825 4048 860 4066
rect 825 4030 834 4048
rect 851 4030 860 4048
rect 825 4012 860 4030
rect 825 3994 834 4012
rect 851 3994 860 4012
rect 825 3976 860 3994
rect 825 3958 834 3976
rect 851 3958 860 3976
rect 825 3940 860 3958
rect 825 3922 834 3940
rect 851 3922 860 3940
rect 825 3904 860 3922
rect 825 3886 834 3904
rect 851 3886 860 3904
rect 825 3868 860 3886
rect 825 3850 834 3868
rect 851 3850 860 3868
rect 825 3832 860 3850
rect 825 3814 834 3832
rect 851 3814 860 3832
rect 825 3796 860 3814
rect 825 3778 834 3796
rect 851 3778 860 3796
rect 825 3760 860 3778
rect 825 3742 834 3760
rect 851 3742 860 3760
rect 825 3724 860 3742
rect 825 3706 834 3724
rect 851 3706 860 3724
rect 825 3688 860 3706
rect 825 3670 834 3688
rect 851 3670 860 3688
rect 825 3652 860 3670
rect 825 3634 834 3652
rect 851 3634 860 3652
rect 825 3616 860 3634
rect 825 3598 834 3616
rect 851 3598 860 3616
rect 825 3580 860 3598
rect 825 3562 834 3580
rect 851 3562 860 3580
rect 825 3544 860 3562
rect 825 3526 834 3544
rect 851 3526 860 3544
rect 825 3508 860 3526
rect 825 3490 834 3508
rect 851 3490 860 3508
rect 825 3472 860 3490
rect 825 3454 834 3472
rect 851 3454 860 3472
rect 825 3436 860 3454
rect 825 3418 834 3436
rect 851 3418 860 3436
rect 825 3400 860 3418
rect 825 3382 834 3400
rect 851 3382 860 3400
rect 825 3364 860 3382
rect 825 3346 834 3364
rect 851 3346 860 3364
rect 825 3328 860 3346
rect 825 3310 834 3328
rect 851 3310 860 3328
rect 825 3292 860 3310
rect 825 3274 834 3292
rect 851 3274 860 3292
rect 825 3256 860 3274
rect 825 3238 834 3256
rect 851 3238 860 3256
rect 825 3220 860 3238
rect 825 3202 834 3220
rect 851 3202 860 3220
rect 825 3184 860 3202
rect 825 3166 834 3184
rect 851 3166 860 3184
rect 825 3148 860 3166
rect 825 3130 834 3148
rect 851 3130 860 3148
rect 825 3112 860 3130
rect 825 3094 834 3112
rect 851 3094 860 3112
rect 825 3076 860 3094
rect 825 3058 834 3076
rect 851 3058 860 3076
rect 825 3040 860 3058
rect 825 3022 834 3040
rect 851 3022 860 3040
rect 825 3004 860 3022
rect 825 2986 834 3004
rect 851 2986 860 3004
rect 825 2968 860 2986
rect 825 2950 834 2968
rect 851 2950 860 2968
rect 825 2932 860 2950
rect 825 2914 834 2932
rect 851 2914 860 2932
rect 825 2896 860 2914
rect 825 2878 834 2896
rect 851 2878 860 2896
rect 825 2860 860 2878
rect 825 2842 834 2860
rect 851 2842 860 2860
rect 825 2824 860 2842
rect 825 2806 834 2824
rect 851 2806 860 2824
rect 825 2788 860 2806
rect 825 2770 834 2788
rect 851 2770 860 2788
rect 825 2752 860 2770
rect 825 2734 834 2752
rect 851 2734 860 2752
rect 825 2716 860 2734
rect 825 2698 834 2716
rect 851 2698 860 2716
rect 825 2680 860 2698
rect 825 2662 834 2680
rect 851 2662 860 2680
rect 825 2644 860 2662
rect 825 2626 834 2644
rect 851 2626 860 2644
rect 825 2608 860 2626
rect 825 2590 834 2608
rect 851 2590 860 2608
rect 825 2572 860 2590
rect 825 2554 834 2572
rect 851 2554 860 2572
rect 825 2536 860 2554
rect 825 2518 834 2536
rect 851 2518 860 2536
rect 825 2500 860 2518
rect 825 2482 834 2500
rect 851 2482 860 2500
rect 825 2464 860 2482
rect 825 2446 834 2464
rect 851 2446 860 2464
rect 825 2428 860 2446
rect 825 2410 834 2428
rect 851 2410 860 2428
rect 825 2392 860 2410
rect 825 2374 834 2392
rect 851 2374 860 2392
rect 825 2356 860 2374
rect 825 2338 834 2356
rect 851 2338 860 2356
rect 825 2320 860 2338
rect 825 2302 834 2320
rect 851 2302 860 2320
rect 825 2284 860 2302
rect 825 2266 834 2284
rect 851 2266 860 2284
rect 825 2248 860 2266
rect 825 2230 834 2248
rect 851 2230 860 2248
rect 825 2212 860 2230
rect 825 2194 834 2212
rect 851 2194 860 2212
rect 825 2176 860 2194
rect 825 2158 834 2176
rect 851 2158 860 2176
rect 825 2140 860 2158
rect 825 2122 834 2140
rect 851 2122 860 2140
rect 825 2104 860 2122
rect 825 2086 834 2104
rect 851 2086 860 2104
rect 825 2068 860 2086
rect 825 2050 834 2068
rect 851 2050 860 2068
rect 825 2032 860 2050
rect 825 2014 834 2032
rect 851 2014 860 2032
rect 825 1996 860 2014
rect 825 1978 834 1996
rect 851 1978 860 1996
rect 825 1960 860 1978
rect 825 1942 834 1960
rect 851 1942 860 1960
rect 825 1924 860 1942
rect 825 1906 834 1924
rect 851 1906 860 1924
rect 825 1888 860 1906
rect 825 1870 834 1888
rect 851 1870 860 1888
rect 825 1852 860 1870
rect 825 1834 834 1852
rect 851 1834 860 1852
rect 825 1816 860 1834
rect 825 1798 834 1816
rect 851 1798 860 1816
rect 825 1780 860 1798
rect 825 1762 834 1780
rect 851 1762 860 1780
rect 825 1744 860 1762
rect 825 1726 834 1744
rect 851 1726 860 1744
rect 825 1708 860 1726
rect 825 1690 834 1708
rect 851 1690 860 1708
rect 825 1672 860 1690
rect 825 1654 834 1672
rect 851 1654 860 1672
rect 825 1636 860 1654
rect 825 1618 834 1636
rect 851 1618 860 1636
rect 825 1600 860 1618
rect 825 1582 834 1600
rect 851 1582 860 1600
rect 825 1564 860 1582
rect 825 1546 834 1564
rect 851 1546 860 1564
rect 825 1528 860 1546
rect 825 1510 834 1528
rect 851 1510 860 1528
rect 825 1492 860 1510
rect 825 1474 834 1492
rect 851 1474 860 1492
rect 825 1456 860 1474
rect 825 1438 834 1456
rect 851 1438 860 1456
rect 825 1420 860 1438
rect 825 1402 834 1420
rect 851 1402 860 1420
rect 825 1384 860 1402
rect 825 1366 834 1384
rect 851 1366 860 1384
rect 825 1348 860 1366
rect 825 1330 834 1348
rect 851 1330 860 1348
rect 825 1312 860 1330
rect 825 1294 834 1312
rect 851 1294 860 1312
rect 825 1276 860 1294
rect 825 1258 834 1276
rect 851 1258 860 1276
rect 825 1240 860 1258
rect 825 1222 834 1240
rect 851 1222 860 1240
rect 825 1204 860 1222
rect 825 1186 834 1204
rect 851 1186 860 1204
rect 825 1168 860 1186
rect 825 1150 834 1168
rect 851 1150 860 1168
rect 825 1132 860 1150
rect 825 1114 834 1132
rect 851 1114 860 1132
rect 825 1096 860 1114
rect 825 1078 834 1096
rect 851 1078 860 1096
rect 825 1060 860 1078
rect 825 1042 834 1060
rect 851 1042 860 1060
rect 825 1024 860 1042
rect 825 1006 834 1024
rect 851 1006 860 1024
rect 825 988 860 1006
rect 825 970 834 988
rect 851 970 860 988
rect 825 952 860 970
rect 825 934 834 952
rect 851 934 860 952
rect 825 916 860 934
rect 825 898 834 916
rect 851 898 860 916
rect 825 880 860 898
rect 825 862 834 880
rect 851 862 860 880
rect 825 844 860 862
rect 825 826 834 844
rect 851 826 860 844
rect 825 808 860 826
rect 825 790 834 808
rect 851 790 860 808
rect 825 772 860 790
rect 825 754 834 772
rect 851 754 860 772
rect 825 736 860 754
rect 825 718 834 736
rect 851 718 860 736
rect 825 700 860 718
rect 825 682 834 700
rect 851 682 860 700
rect 825 664 860 682
rect 825 646 834 664
rect 851 646 860 664
rect 825 628 860 646
rect 825 610 834 628
rect 851 610 860 628
rect 825 601 860 610
<< mvndiffc >>
rect 199 4750 216 4768
rect 199 4714 216 4732
rect 199 4678 216 4696
rect 199 4642 216 4660
rect 199 4606 216 4624
rect 199 4570 216 4588
rect 199 4534 216 4552
rect 199 4498 216 4516
rect 199 4462 216 4480
rect 199 4426 216 4444
rect 199 4390 216 4408
rect 199 4354 216 4372
rect 199 4318 216 4336
rect 199 4282 216 4300
rect 199 4246 216 4264
rect 199 4210 216 4228
rect 199 4174 216 4192
rect 199 4138 216 4156
rect 199 4102 216 4120
rect 199 4066 216 4084
rect 199 4030 216 4048
rect 199 3994 216 4012
rect 199 3958 216 3976
rect 199 3922 216 3940
rect 199 3886 216 3904
rect 199 3850 216 3868
rect 199 3814 216 3832
rect 199 3778 216 3796
rect 199 3742 216 3760
rect 199 3706 216 3724
rect 199 3670 216 3688
rect 199 3634 216 3652
rect 199 3598 216 3616
rect 199 3562 216 3580
rect 199 3526 216 3544
rect 199 3490 216 3508
rect 199 3454 216 3472
rect 199 3418 216 3436
rect 199 3382 216 3400
rect 199 3346 216 3364
rect 199 3310 216 3328
rect 199 3274 216 3292
rect 199 3238 216 3256
rect 199 3202 216 3220
rect 199 3166 216 3184
rect 199 3130 216 3148
rect 199 3094 216 3112
rect 199 3058 216 3076
rect 199 3022 216 3040
rect 199 2986 216 3004
rect 199 2950 216 2968
rect 199 2914 216 2932
rect 199 2878 216 2896
rect 199 2842 216 2860
rect 199 2806 216 2824
rect 199 2770 216 2788
rect 199 2734 216 2752
rect 199 2698 216 2716
rect 199 2662 216 2680
rect 199 2626 216 2644
rect 199 2590 216 2608
rect 199 2554 216 2572
rect 199 2518 216 2536
rect 199 2482 216 2500
rect 199 2446 216 2464
rect 199 2410 216 2428
rect 199 2374 216 2392
rect 199 2338 216 2356
rect 199 2302 216 2320
rect 199 2266 216 2284
rect 199 2230 216 2248
rect 199 2194 216 2212
rect 199 2158 216 2176
rect 199 2122 216 2140
rect 199 2086 216 2104
rect 199 2050 216 2068
rect 199 2014 216 2032
rect 199 1978 216 1996
rect 199 1942 216 1960
rect 199 1906 216 1924
rect 199 1870 216 1888
rect 199 1834 216 1852
rect 199 1798 216 1816
rect 199 1762 216 1780
rect 199 1726 216 1744
rect 199 1690 216 1708
rect 199 1654 216 1672
rect 199 1618 216 1636
rect 199 1582 216 1600
rect 199 1546 216 1564
rect 199 1510 216 1528
rect 199 1474 216 1492
rect 199 1438 216 1456
rect 199 1402 216 1420
rect 199 1366 216 1384
rect 199 1330 216 1348
rect 199 1294 216 1312
rect 199 1258 216 1276
rect 199 1222 216 1240
rect 199 1186 216 1204
rect 199 1150 216 1168
rect 199 1114 216 1132
rect 199 1078 216 1096
rect 199 1042 216 1060
rect 199 1006 216 1024
rect 199 970 216 988
rect 199 934 216 952
rect 199 898 216 916
rect 199 862 216 880
rect 199 826 216 844
rect 199 790 216 808
rect 199 754 216 772
rect 199 718 216 736
rect 199 682 216 700
rect 199 646 216 664
rect 199 610 216 628
rect 834 4750 851 4768
rect 834 4714 851 4732
rect 834 4678 851 4696
rect 834 4642 851 4660
rect 834 4606 851 4624
rect 834 4570 851 4588
rect 834 4534 851 4552
rect 834 4498 851 4516
rect 834 4462 851 4480
rect 834 4426 851 4444
rect 834 4390 851 4408
rect 834 4354 851 4372
rect 834 4318 851 4336
rect 834 4282 851 4300
rect 834 4246 851 4264
rect 834 4210 851 4228
rect 834 4174 851 4192
rect 834 4138 851 4156
rect 834 4102 851 4120
rect 834 4066 851 4084
rect 834 4030 851 4048
rect 834 3994 851 4012
rect 834 3958 851 3976
rect 834 3922 851 3940
rect 834 3886 851 3904
rect 834 3850 851 3868
rect 834 3814 851 3832
rect 834 3778 851 3796
rect 834 3742 851 3760
rect 834 3706 851 3724
rect 834 3670 851 3688
rect 834 3634 851 3652
rect 834 3598 851 3616
rect 834 3562 851 3580
rect 834 3526 851 3544
rect 834 3490 851 3508
rect 834 3454 851 3472
rect 834 3418 851 3436
rect 834 3382 851 3400
rect 834 3346 851 3364
rect 834 3310 851 3328
rect 834 3274 851 3292
rect 834 3238 851 3256
rect 834 3202 851 3220
rect 834 3166 851 3184
rect 834 3130 851 3148
rect 834 3094 851 3112
rect 834 3058 851 3076
rect 834 3022 851 3040
rect 834 2986 851 3004
rect 834 2950 851 2968
rect 834 2914 851 2932
rect 834 2878 851 2896
rect 834 2842 851 2860
rect 834 2806 851 2824
rect 834 2770 851 2788
rect 834 2734 851 2752
rect 834 2698 851 2716
rect 834 2662 851 2680
rect 834 2626 851 2644
rect 834 2590 851 2608
rect 834 2554 851 2572
rect 834 2518 851 2536
rect 834 2482 851 2500
rect 834 2446 851 2464
rect 834 2410 851 2428
rect 834 2374 851 2392
rect 834 2338 851 2356
rect 834 2302 851 2320
rect 834 2266 851 2284
rect 834 2230 851 2248
rect 834 2194 851 2212
rect 834 2158 851 2176
rect 834 2122 851 2140
rect 834 2086 851 2104
rect 834 2050 851 2068
rect 834 2014 851 2032
rect 834 1978 851 1996
rect 834 1942 851 1960
rect 834 1906 851 1924
rect 834 1870 851 1888
rect 834 1834 851 1852
rect 834 1798 851 1816
rect 834 1762 851 1780
rect 834 1726 851 1744
rect 834 1690 851 1708
rect 834 1654 851 1672
rect 834 1618 851 1636
rect 834 1582 851 1600
rect 834 1546 851 1564
rect 834 1510 851 1528
rect 834 1474 851 1492
rect 834 1438 851 1456
rect 834 1402 851 1420
rect 834 1366 851 1384
rect 834 1330 851 1348
rect 834 1294 851 1312
rect 834 1258 851 1276
rect 834 1222 851 1240
rect 834 1186 851 1204
rect 834 1150 851 1168
rect 834 1114 851 1132
rect 834 1078 851 1096
rect 834 1042 851 1060
rect 834 1006 851 1024
rect 834 970 851 988
rect 834 934 851 952
rect 834 898 851 916
rect 834 862 851 880
rect 834 826 851 844
rect 834 790 851 808
rect 834 754 851 772
rect 834 718 851 736
rect 834 682 851 700
rect 834 646 851 664
rect 834 610 851 628
<< poly >>
rect 225 4801 825 4852
rect 225 550 825 601
<< locali >>
rect 199 4768 216 4801
rect 199 4732 216 4750
rect 199 4696 216 4714
rect 199 4660 216 4678
rect 199 4624 216 4642
rect 199 4588 216 4606
rect 199 4552 216 4570
rect 199 4516 216 4534
rect 199 4480 216 4498
rect 199 4444 216 4462
rect 199 4408 216 4426
rect 199 4372 216 4390
rect 199 4336 216 4354
rect 199 4300 216 4318
rect 199 4264 216 4282
rect 199 4228 216 4246
rect 199 4192 216 4210
rect 199 4156 216 4174
rect 199 4120 216 4138
rect 199 4084 216 4102
rect 199 4048 216 4066
rect 199 4012 216 4030
rect 199 3976 216 3994
rect 199 3940 216 3958
rect 199 3904 216 3922
rect 199 3868 216 3886
rect 199 3832 216 3850
rect 199 3796 216 3814
rect 199 3760 216 3778
rect 199 3724 216 3742
rect 199 3688 216 3706
rect 199 3652 216 3670
rect 199 3616 216 3634
rect 199 3580 216 3598
rect 199 3544 216 3562
rect 199 3508 216 3526
rect 199 3472 216 3490
rect 199 3436 216 3454
rect 199 3400 216 3418
rect 199 3364 216 3382
rect 199 3328 216 3346
rect 199 3292 216 3310
rect 199 3256 216 3274
rect 199 3220 216 3238
rect 199 3184 216 3202
rect 199 3148 216 3166
rect 199 3112 216 3130
rect 199 3076 216 3094
rect 199 3040 216 3058
rect 199 3004 216 3022
rect 199 2968 216 2986
rect 199 2932 216 2950
rect 199 2896 216 2914
rect 199 2860 216 2878
rect 199 2824 216 2842
rect 199 2788 216 2806
rect 199 2752 216 2770
rect 199 2716 216 2734
rect 199 2680 216 2698
rect 199 2644 216 2662
rect 199 2608 216 2626
rect 199 2572 216 2590
rect 199 2536 216 2554
rect 199 2500 216 2518
rect 199 2464 216 2482
rect 199 2428 216 2446
rect 199 2392 216 2410
rect 199 2356 216 2374
rect 199 2320 216 2338
rect 199 2284 216 2302
rect 199 2248 216 2266
rect 199 2212 216 2230
rect 199 2176 216 2194
rect 199 2140 216 2158
rect 199 2104 216 2122
rect 199 2068 216 2086
rect 199 2032 216 2050
rect 199 1996 216 2014
rect 199 1960 216 1978
rect 199 1924 216 1942
rect 199 1888 216 1906
rect 199 1852 216 1870
rect 199 1816 216 1834
rect 199 1780 216 1798
rect 199 1744 216 1762
rect 199 1708 216 1726
rect 199 1672 216 1690
rect 199 1636 216 1654
rect 199 1600 216 1618
rect 199 1564 216 1582
rect 199 1528 216 1546
rect 199 1492 216 1510
rect 199 1456 216 1474
rect 199 1420 216 1438
rect 199 1384 216 1402
rect 199 1348 216 1366
rect 199 1312 216 1330
rect 199 1276 216 1294
rect 199 1240 216 1258
rect 199 1204 216 1222
rect 199 1168 216 1186
rect 199 1132 216 1150
rect 199 1096 216 1114
rect 199 1060 216 1078
rect 199 1024 216 1042
rect 199 988 216 1006
rect 199 952 216 970
rect 199 916 216 934
rect 199 880 216 898
rect 199 844 216 862
rect 199 808 216 826
rect 199 772 216 790
rect 199 736 216 754
rect 199 700 216 718
rect 199 664 216 682
rect 199 628 216 646
rect 199 601 216 610
rect 834 4768 851 4801
rect 834 4732 851 4750
rect 834 4696 851 4714
rect 834 4660 851 4678
rect 834 4624 851 4642
rect 834 4588 851 4606
rect 834 4552 851 4570
rect 834 4516 851 4534
rect 834 4480 851 4498
rect 834 4444 851 4462
rect 834 4408 851 4426
rect 834 4372 851 4390
rect 834 4336 851 4354
rect 834 4300 851 4318
rect 834 4264 851 4282
rect 834 4228 851 4246
rect 834 4192 851 4210
rect 834 4156 851 4174
rect 834 4120 851 4138
rect 834 4084 851 4102
rect 834 4048 851 4066
rect 834 4012 851 4030
rect 834 3976 851 3994
rect 834 3940 851 3958
rect 834 3904 851 3922
rect 834 3868 851 3886
rect 834 3832 851 3850
rect 834 3796 851 3814
rect 834 3760 851 3778
rect 834 3724 851 3742
rect 834 3688 851 3706
rect 834 3652 851 3670
rect 834 3616 851 3634
rect 834 3580 851 3598
rect 834 3544 851 3562
rect 834 3508 851 3526
rect 834 3472 851 3490
rect 834 3436 851 3454
rect 834 3400 851 3418
rect 834 3364 851 3382
rect 834 3328 851 3346
rect 834 3292 851 3310
rect 834 3256 851 3274
rect 834 3220 851 3238
rect 834 3184 851 3202
rect 834 3148 851 3166
rect 834 3112 851 3130
rect 834 3076 851 3094
rect 834 3040 851 3058
rect 834 3004 851 3022
rect 834 2968 851 2986
rect 834 2932 851 2950
rect 834 2896 851 2914
rect 834 2860 851 2878
rect 834 2824 851 2842
rect 834 2788 851 2806
rect 834 2752 851 2770
rect 834 2716 851 2734
rect 834 2680 851 2698
rect 834 2644 851 2662
rect 834 2608 851 2626
rect 834 2572 851 2590
rect 834 2536 851 2554
rect 834 2500 851 2518
rect 834 2464 851 2482
rect 834 2428 851 2446
rect 834 2392 851 2410
rect 834 2356 851 2374
rect 834 2320 851 2338
rect 834 2284 851 2302
rect 834 2248 851 2266
rect 834 2212 851 2230
rect 834 2176 851 2194
rect 834 2140 851 2158
rect 834 2104 851 2122
rect 834 2068 851 2086
rect 834 2032 851 2050
rect 834 1996 851 2014
rect 834 1960 851 1978
rect 834 1924 851 1942
rect 834 1888 851 1906
rect 834 1852 851 1870
rect 834 1816 851 1834
rect 834 1780 851 1798
rect 834 1744 851 1762
rect 834 1708 851 1726
rect 834 1672 851 1690
rect 834 1636 851 1654
rect 834 1600 851 1618
rect 834 1564 851 1582
rect 834 1528 851 1546
rect 834 1492 851 1510
rect 834 1456 851 1474
rect 834 1420 851 1438
rect 834 1384 851 1402
rect 834 1348 851 1366
rect 834 1312 851 1330
rect 834 1276 851 1294
rect 834 1240 851 1258
rect 834 1204 851 1222
rect 834 1168 851 1186
rect 834 1132 851 1150
rect 834 1096 851 1114
rect 834 1060 851 1078
rect 834 1024 851 1042
rect 834 988 851 1006
rect 834 952 851 970
rect 834 916 851 934
rect 834 880 851 898
rect 834 844 851 862
rect 834 808 851 826
rect 834 772 851 790
rect 834 736 851 754
rect 834 700 851 718
rect 834 664 851 682
rect 834 628 851 646
rect 834 601 851 610
<< end >>
