magic
tech sky130A
magscale 1 2
timestamp 1621849157
<< nwell >>
rect 0 14540 7636 14770
rect 38 12728 344 14540
rect 2136 13598 6460 14540
rect 2386 13544 6460 13598
rect 2136 10390 6460 13544
<< mvpsubdiff >>
rect 0 -18 100 16
rect 134 -18 300 16
rect 334 -18 500 16
rect 534 -18 700 16
rect 734 -18 900 16
rect 934 -18 1100 16
rect 1134 -18 1300 16
rect 1334 -18 1500 16
rect 1534 -18 1700 16
rect 1734 -18 1900 16
rect 1934 -18 2100 16
rect 2134 -18 2300 16
rect 2334 -18 2500 16
rect 2534 -18 2700 16
rect 2734 -18 2900 16
rect 2934 -18 3100 16
rect 3134 -18 3300 16
rect 3334 -18 3500 16
rect 3534 -18 3700 16
rect 3734 -18 3900 16
rect 3934 -18 4100 16
rect 4134 -18 4300 16
rect 4334 -18 4500 16
rect 4534 -18 4700 16
rect 4734 -18 4900 16
rect 4934 -18 5100 16
rect 5134 -18 5300 16
rect 5334 -18 5500 16
rect 5534 -18 5700 16
rect 5734 -18 5900 16
rect 5934 -18 6100 16
rect 6134 -18 6300 16
rect 6334 -18 6500 16
rect 6534 -18 6700 16
rect 6734 -18 6900 16
rect 6934 -18 7100 16
rect 7134 -18 7300 16
rect 7334 -18 7500 16
rect 7534 -18 7636 16
<< mvnsubdiff >>
rect 66 14670 100 14704
rect 134 14670 300 14704
rect 334 14670 500 14704
rect 534 14670 700 14704
rect 734 14670 900 14704
rect 934 14670 1100 14704
rect 1134 14670 1300 14704
rect 1334 14670 1500 14704
rect 1534 14670 1700 14704
rect 1734 14670 1900 14704
rect 1934 14670 2100 14704
rect 2134 14670 2300 14704
rect 2334 14670 2500 14704
rect 2534 14670 2700 14704
rect 2734 14670 2900 14704
rect 2934 14670 3100 14704
rect 3134 14670 3300 14704
rect 3334 14670 3500 14704
rect 3534 14670 3700 14704
rect 3734 14670 3900 14704
rect 3934 14670 4100 14704
rect 4134 14670 4300 14704
rect 4334 14670 4500 14704
rect 4534 14670 4700 14704
rect 4734 14670 4900 14704
rect 4934 14670 5100 14704
rect 5134 14670 5300 14704
rect 5334 14670 5500 14704
rect 5534 14670 5700 14704
rect 5734 14670 5900 14704
rect 5934 14670 6100 14704
rect 6134 14670 6300 14704
rect 6334 14670 6500 14704
rect 6534 14670 6700 14704
rect 6734 14670 6900 14704
rect 6934 14670 7100 14704
rect 7134 14670 7300 14704
rect 7334 14670 7570 14704
<< mvpsubdiffcont >>
rect 100 -18 134 16
rect 300 -18 334 16
rect 500 -18 534 16
rect 700 -18 734 16
rect 900 -18 934 16
rect 1100 -18 1134 16
rect 1300 -18 1334 16
rect 1500 -18 1534 16
rect 1700 -18 1734 16
rect 1900 -18 1934 16
rect 2100 -18 2134 16
rect 2300 -18 2334 16
rect 2500 -18 2534 16
rect 2700 -18 2734 16
rect 2900 -18 2934 16
rect 3100 -18 3134 16
rect 3300 -18 3334 16
rect 3500 -18 3534 16
rect 3700 -18 3734 16
rect 3900 -18 3934 16
rect 4100 -18 4134 16
rect 4300 -18 4334 16
rect 4500 -18 4534 16
rect 4700 -18 4734 16
rect 4900 -18 4934 16
rect 5100 -18 5134 16
rect 5300 -18 5334 16
rect 5500 -18 5534 16
rect 5700 -18 5734 16
rect 5900 -18 5934 16
rect 6100 -18 6134 16
rect 6300 -18 6334 16
rect 6500 -18 6534 16
rect 6700 -18 6734 16
rect 6900 -18 6934 16
rect 7100 -18 7134 16
rect 7300 -18 7334 16
rect 7500 -18 7534 16
<< mvnsubdiffcont >>
rect 100 14670 134 14704
rect 300 14670 334 14704
rect 500 14670 534 14704
rect 700 14670 734 14704
rect 900 14670 934 14704
rect 1100 14670 1134 14704
rect 1300 14670 1334 14704
rect 1500 14670 1534 14704
rect 1700 14670 1734 14704
rect 1900 14670 1934 14704
rect 2100 14670 2134 14704
rect 2300 14670 2334 14704
rect 2500 14670 2534 14704
rect 2700 14670 2734 14704
rect 2900 14670 2934 14704
rect 3100 14670 3134 14704
rect 3300 14670 3334 14704
rect 3500 14670 3534 14704
rect 3700 14670 3734 14704
rect 3900 14670 3934 14704
rect 4100 14670 4134 14704
rect 4300 14670 4334 14704
rect 4500 14670 4534 14704
rect 4700 14670 4734 14704
rect 4900 14670 4934 14704
rect 5100 14670 5134 14704
rect 5300 14670 5334 14704
rect 5500 14670 5534 14704
rect 5700 14670 5734 14704
rect 5900 14670 5934 14704
rect 6100 14670 6134 14704
rect 6300 14670 6334 14704
rect 6500 14670 6534 14704
rect 6700 14670 6734 14704
rect 6900 14670 6934 14704
rect 7100 14670 7134 14704
rect 7300 14670 7334 14704
<< poly >>
rect 3272 13944 3798 14510
rect 3272 13910 3504 13944
rect 3554 13910 3798 13944
rect 3272 13570 3798 13910
rect 3272 13520 3746 13570
rect 3780 13520 3798 13570
rect 3272 13510 3798 13520
rect 4798 13510 5324 14510
rect 3272 9614 3798 10180
rect 3272 9580 3496 9614
rect 3546 9580 3798 9614
rect 3272 9180 3798 9580
rect 3272 4880 3798 5880
rect 4798 4880 5324 5880
<< polycont >>
rect 3504 13910 3554 13944
rect 3746 13520 3780 13570
rect 1702 10408 1770 10442
rect 3496 9580 3546 9614
rect 2292 9294 2342 9328
rect 1128 9018 1328 9052
rect 6236 5344 6286 5378
rect 290 642 324 692
<< xpolycontact >>
rect 6960 10914 7030 11346
rect 6642 4562 6712 4994
rect 6642 2380 6712 2812
rect 6960 2380 7030 2812
rect 7278 10914 7348 11346
rect 7278 2380 7348 2812
<< xpolyres >>
rect 6642 2812 6712 4562
rect 6960 2812 7030 10914
rect 7278 2812 7348 10914
<< locali >>
rect 0 14670 100 14704
rect 134 14670 300 14704
rect 334 14670 500 14704
rect 534 14670 700 14704
rect 734 14670 900 14704
rect 934 14670 1100 14704
rect 1134 14670 1300 14704
rect 1334 14670 1500 14704
rect 1534 14670 1700 14704
rect 1734 14670 1900 14704
rect 1934 14670 2100 14704
rect 2134 14670 2300 14704
rect 2334 14670 2500 14704
rect 2534 14670 2700 14704
rect 2734 14670 2900 14704
rect 2934 14670 3100 14704
rect 3134 14670 3300 14704
rect 3334 14670 3500 14704
rect 3534 14670 3700 14704
rect 3734 14670 3900 14704
rect 3934 14670 4100 14704
rect 4134 14670 4300 14704
rect 4334 14670 4500 14704
rect 4534 14670 4700 14704
rect 4734 14670 4900 14704
rect 4934 14670 5100 14704
rect 5134 14670 5300 14704
rect 5334 14670 5500 14704
rect 5534 14670 5700 14704
rect 5734 14670 5900 14704
rect 5934 14670 6100 14704
rect 6134 14670 6300 14704
rect 6334 14670 6500 14704
rect 6534 14670 6700 14704
rect 6734 14670 6900 14704
rect 6934 14670 7100 14704
rect 7134 14670 7300 14704
rect 7334 14670 7500 14704
rect 7534 14670 7636 14704
rect 174 12648 208 14670
rect 1584 13910 3144 13944
rect 3194 13910 3210 13944
rect 1584 11092 1618 13910
rect 3290 13460 3324 14670
rect 3380 13910 3396 13944
rect 3446 13910 3504 13944
rect 3554 13910 3578 13944
rect 3746 13570 3780 13586
rect 3746 13460 3780 13520
rect 4816 13460 4850 14670
rect 6342 13460 6376 14670
rect 6958 11346 7032 11348
rect 6958 10914 6960 11346
rect 7030 11144 7032 11346
rect 7276 11346 7350 11348
rect 7276 11144 7278 11346
rect 7030 11110 7278 11144
rect 7030 10914 7032 11110
rect 6958 10912 7032 10914
rect 7276 10914 7278 11110
rect 7348 10914 7350 11346
rect 7276 10912 7350 10914
rect 1854 10444 1888 10492
rect 412 10408 1702 10442
rect 1770 10408 1786 10442
rect 1854 10410 2034 10444
rect 290 692 324 708
rect 174 494 208 544
rect 290 494 324 642
rect 412 494 446 10408
rect 2000 9914 2034 10410
rect 2220 10436 2254 10460
rect 2220 10380 2254 10386
rect 3746 10436 3780 10460
rect 3746 10380 3780 10386
rect 5272 10436 5306 10460
rect 5272 10380 5306 10386
rect 2000 9852 2034 9864
rect 1216 9580 3496 9614
rect 3546 9580 3562 9614
rect 1216 9052 1250 9580
rect 2220 9294 2292 9328
rect 2342 9294 2358 9328
rect 2000 9250 2034 9258
rect 1112 9018 1128 9052
rect 1328 9018 1344 9052
rect 584 494 618 562
rect 174 460 618 494
rect 1854 494 1888 562
rect 2000 494 2034 9200
rect 2220 9202 2254 9294
rect 2220 9130 2254 9152
rect 3746 9202 3780 9290
rect 3746 9130 3780 9152
rect 3290 6106 3324 6130
rect 3290 6050 3324 6056
rect 4816 6106 4850 6130
rect 4816 6050 4850 6056
rect 6220 5344 6236 5378
rect 6286 5344 6324 5378
rect 3746 4996 6714 5030
rect 3290 4904 3324 4910
rect 3290 4830 3324 4854
rect 3746 4830 3780 4996
rect 6640 4994 6714 4996
rect 4816 4904 4850 4910
rect 4816 4830 4850 4854
rect 5272 4904 5306 4910
rect 5272 4830 5306 4854
rect 6640 4562 6642 4994
rect 6712 4562 6714 4994
rect 6640 4560 6714 4562
rect 6640 2812 6714 2814
rect 2220 2406 2254 2430
rect 2220 2350 2254 2356
rect 6342 2362 6376 2430
rect 6342 2300 6376 2312
rect 6640 2380 6642 2812
rect 6712 2380 6714 2812
rect 6640 2272 6714 2380
rect 6958 2812 7032 2814
rect 6958 2380 6960 2812
rect 7030 2380 7032 2812
rect 6958 2362 7032 2380
rect 6958 2312 6978 2362
rect 7012 2312 7032 2362
rect 6958 2300 7032 2312
rect 7276 2812 7350 2814
rect 7276 2380 7278 2812
rect 7348 2380 7350 2812
rect 7276 2360 7350 2380
rect 7276 2310 7296 2360
rect 7330 2310 7350 2360
rect 7276 2300 7350 2310
rect 6640 2222 6660 2272
rect 6694 2222 6714 2272
rect 6640 2212 6714 2222
rect 2538 1376 2610 1440
rect 3336 1376 3408 1440
rect 4134 1376 4206 1440
rect 4932 1376 5004 1440
rect 5730 1376 5802 1440
rect 2202 1260 6138 1276
rect 2202 1226 6286 1260
rect 2202 1204 6138 1226
rect 2538 560 2610 624
rect 3336 560 3408 624
rect 4134 560 4206 624
rect 4932 560 5004 624
rect 5730 560 5802 624
rect 1854 460 2034 494
rect 2000 16 2034 460
rect 6252 16 6286 1226
rect 0 -18 100 16
rect 134 -18 300 16
rect 334 -18 500 16
rect 534 -18 700 16
rect 734 -18 900 16
rect 934 -18 1100 16
rect 1134 -18 1300 16
rect 1334 -18 1500 16
rect 1534 -18 1700 16
rect 1734 -18 1900 16
rect 1934 -18 2100 16
rect 2134 -18 2300 16
rect 2334 -18 2500 16
rect 2534 -18 2700 16
rect 2734 -18 2900 16
rect 2934 -18 3100 16
rect 3134 -18 3300 16
rect 3334 -18 3500 16
rect 3534 -18 3700 16
rect 3734 -18 3900 16
rect 3934 -18 4100 16
rect 4134 -18 4300 16
rect 4334 -18 4500 16
rect 4534 -18 4700 16
rect 4734 -18 4900 16
rect 4934 -18 5100 16
rect 5134 -18 5300 16
rect 5334 -18 5500 16
rect 5534 -18 5700 16
rect 5734 -18 5900 16
rect 5934 -18 6100 16
rect 6134 -18 6300 16
rect 6334 -18 6500 16
rect 6534 -18 6700 16
rect 6734 -18 6900 16
rect 6934 -18 7100 16
rect 7134 -18 7300 16
rect 7334 -18 7500 16
rect 7534 -18 7636 16
<< viali >>
rect 100 14670 134 14704
rect 300 14670 334 14704
rect 500 14670 534 14704
rect 700 14670 734 14704
rect 900 14670 934 14704
rect 1100 14670 1134 14704
rect 1300 14670 1334 14704
rect 1500 14670 1534 14704
rect 1700 14670 1734 14704
rect 1900 14670 1934 14704
rect 2100 14670 2134 14704
rect 2300 14670 2334 14704
rect 2500 14670 2534 14704
rect 2700 14670 2734 14704
rect 2900 14670 2934 14704
rect 3100 14670 3134 14704
rect 3300 14670 3334 14704
rect 3500 14670 3534 14704
rect 3700 14670 3734 14704
rect 3900 14670 3934 14704
rect 4100 14670 4134 14704
rect 4300 14670 4334 14704
rect 4500 14670 4534 14704
rect 4700 14670 4734 14704
rect 4900 14670 4934 14704
rect 5100 14670 5134 14704
rect 5300 14670 5334 14704
rect 5500 14670 5534 14704
rect 5700 14670 5734 14704
rect 5900 14670 5934 14704
rect 6100 14670 6134 14704
rect 6300 14670 6334 14704
rect 6500 14670 6534 14704
rect 6700 14670 6734 14704
rect 6900 14670 6934 14704
rect 7100 14670 7134 14704
rect 7300 14670 7334 14704
rect 7500 14670 7534 14704
rect 3144 13910 3194 13944
rect 3396 13910 3446 13944
rect 2220 10386 2254 10436
rect 3746 10386 3780 10436
rect 5272 10386 5306 10436
rect 2000 9864 2034 9914
rect 2000 9200 2034 9250
rect 2220 9152 2254 9202
rect 3746 9152 3780 9202
rect 3290 6056 3324 6106
rect 4816 6056 4850 6106
rect 3290 4854 3324 4904
rect 4816 4854 4850 4904
rect 5272 4854 5306 4904
rect 2220 2356 2254 2406
rect 6342 2312 6376 2362
rect 6978 2312 7012 2362
rect 7296 2310 7330 2360
rect 6660 2222 6694 2272
rect 100 -18 134 16
rect 300 -18 334 16
rect 500 -18 534 16
rect 700 -18 734 16
rect 900 -18 934 16
rect 1100 -18 1134 16
rect 1300 -18 1334 16
rect 1500 -18 1534 16
rect 1700 -18 1734 16
rect 1900 -18 1934 16
rect 2100 -18 2134 16
rect 2300 -18 2334 16
rect 2500 -18 2534 16
rect 2700 -18 2734 16
rect 2900 -18 2934 16
rect 3100 -18 3134 16
rect 3300 -18 3334 16
rect 3500 -18 3534 16
rect 3700 -18 3734 16
rect 3900 -18 3934 16
rect 4100 -18 4134 16
rect 4300 -18 4334 16
rect 4500 -18 4534 16
rect 4700 -18 4734 16
rect 4900 -18 4934 16
rect 5100 -18 5134 16
rect 5300 -18 5334 16
rect 5500 -18 5534 16
rect 5700 -18 5734 16
rect 5900 -18 5934 16
rect 6100 -18 6134 16
rect 6300 -18 6334 16
rect 6500 -18 6534 16
rect 6700 -18 6734 16
rect 6900 -18 6934 16
rect 7100 -18 7134 16
rect 7300 -18 7334 16
rect 7500 -18 7534 16
<< metal1 >>
rect 0 14704 7636 14736
rect 0 14670 100 14704
rect 134 14670 300 14704
rect 334 14670 500 14704
rect 534 14670 700 14704
rect 734 14670 900 14704
rect 934 14670 1100 14704
rect 1134 14670 1300 14704
rect 1334 14670 1500 14704
rect 1534 14670 1700 14704
rect 1734 14670 1900 14704
rect 1934 14670 2100 14704
rect 2134 14670 2300 14704
rect 2334 14670 2500 14704
rect 2534 14670 2700 14704
rect 2734 14670 2900 14704
rect 2934 14670 3100 14704
rect 3134 14670 3300 14704
rect 3334 14670 3500 14704
rect 3534 14670 3700 14704
rect 3734 14670 3900 14704
rect 3934 14670 4100 14704
rect 4134 14670 4300 14704
rect 4334 14670 4500 14704
rect 4534 14670 4700 14704
rect 4734 14670 4900 14704
rect 4934 14670 5100 14704
rect 5134 14670 5300 14704
rect 5334 14670 5500 14704
rect 5534 14670 5700 14704
rect 5734 14670 5900 14704
rect 5934 14670 6100 14704
rect 6134 14670 6300 14704
rect 6334 14670 6500 14704
rect 6534 14670 6700 14704
rect 6734 14670 6900 14704
rect 6934 14670 7100 14704
rect 7134 14670 7300 14704
rect 7334 14670 7500 14704
rect 7534 14670 7636 14704
rect 0 14640 7636 14670
rect 3100 13944 3458 13958
rect 3100 13910 3144 13944
rect 3194 13910 3396 13944
rect 3446 13910 3458 13944
rect 3100 13898 3458 13910
rect 2206 10436 2266 10450
rect 2206 10386 2220 10436
rect 2254 10386 2266 10436
rect 1988 9914 2048 9928
rect 1988 9864 2000 9914
rect 2034 9864 2048 9914
rect 1988 9250 2048 9864
rect 1988 9200 2000 9250
rect 2034 9200 2048 9250
rect 1988 9186 2048 9200
rect 2206 9202 2266 10386
rect 2206 9152 2220 9202
rect 2254 9152 2266 9202
rect 2206 9140 2266 9152
rect 3732 10436 3792 10450
rect 3732 10386 3746 10436
rect 3780 10386 3792 10436
rect 3732 9202 3792 10386
rect 3732 9152 3746 9202
rect 3780 9152 3792 9202
rect 3732 9140 3792 9152
rect 5258 10436 5318 10450
rect 5258 10386 5272 10436
rect 5306 10386 5318 10436
rect 3278 6106 3338 6120
rect 3278 6056 3290 6106
rect 3324 6056 3338 6106
rect 3278 4904 3338 6056
rect 3278 4854 3290 4904
rect 3324 4854 3338 4904
rect 3278 4840 3338 4854
rect 4804 6106 4864 6120
rect 4804 6056 4816 6106
rect 4850 6056 4864 6106
rect 4804 4904 4864 6056
rect 4804 4854 4816 4904
rect 4850 4854 4864 4904
rect 4804 4840 4864 4854
rect 5258 4904 5318 10386
rect 5258 4854 5272 4904
rect 5306 4854 5318 4904
rect 5258 4840 5318 4854
rect 2206 2406 2266 2420
rect 2206 2356 2220 2406
rect 2254 2356 2266 2406
rect 2206 2226 2266 2356
rect 6330 2362 7024 2368
rect 6330 2312 6342 2362
rect 6376 2312 6978 2362
rect 7012 2312 7024 2362
rect 6330 2306 7024 2312
rect 7282 2360 7342 2372
rect 7282 2310 7296 2360
rect 7330 2310 7342 2360
rect 4140 2272 6714 2278
rect 2206 2166 2604 2226
rect 2544 1730 2604 2166
rect 4140 2222 6660 2272
rect 6694 2222 6714 2272
rect 4140 2216 6714 2222
rect 4140 2130 4200 2216
rect 2916 2070 5796 2130
rect 2916 862 2976 2070
rect 3342 1730 3402 2070
rect 3714 862 3774 2070
rect 4140 1730 4200 2070
rect 4512 862 4572 2070
rect 4938 1730 4998 2070
rect 5310 862 5370 2070
rect 5736 1730 5796 2070
rect 7282 862 7342 2310
rect 2656 802 2976 862
rect 3454 802 3774 862
rect 4252 802 4572 862
rect 5050 802 5370 862
rect 5848 802 7342 862
rect 0 16 7636 48
rect 0 -18 100 16
rect 134 -18 300 16
rect 334 -18 500 16
rect 534 -18 700 16
rect 734 -18 900 16
rect 934 -18 1100 16
rect 1134 -18 1300 16
rect 1334 -18 1500 16
rect 1534 -18 1700 16
rect 1734 -18 1900 16
rect 1934 -18 2100 16
rect 2134 -18 2300 16
rect 2334 -18 2500 16
rect 2534 -18 2700 16
rect 2734 -18 2900 16
rect 2934 -18 3100 16
rect 3134 -18 3300 16
rect 3334 -18 3500 16
rect 3534 -18 3700 16
rect 3734 -18 3900 16
rect 3934 -18 4100 16
rect 4134 -18 4300 16
rect 4334 -18 4500 16
rect 4534 -18 4700 16
rect 4734 -18 4900 16
rect 4934 -18 5100 16
rect 5134 -18 5300 16
rect 5334 -18 5500 16
rect 5534 -18 5700 16
rect 5734 -18 5900 16
rect 5934 -18 6100 16
rect 6134 -18 6300 16
rect 6334 -18 6500 16
rect 6534 -18 6700 16
rect 6734 -18 6900 16
rect 6934 -18 7100 16
rect 7134 -18 7300 16
rect 7334 -18 7500 16
rect 7534 -18 7636 16
rect 0 -48 7636 -18
use sc_pmos  sc_pmos_0
timestamp 1616540248
transform 1 0 -360 0 1 -2468
box 400 2928 700 15200
use sc_nmos_426  sc_nmos_426_0
timestamp 1616700505
transform 1 0 186 0 1 -640
box 380 1100 1720 9704
use sc_nmos_31  sc_nmos_31_0
timestamp 1616174596
transform 1 0 1186 0 1 9290
box 380 1100 720 1904
use sky130_fd_pr__pnp_05v5_W3p40L3p40  sky130_fd_pr__pnp_05v5_W3p40L3p40_0
timestamp 1615375237
transform 1 0 2176 0 1 1250
box 26 26 770 795
use sky130_fd_pr__pnp_05v5_W3p40L3p40  sky130_fd_pr__pnp_05v5_W3p40L3p40_2
timestamp 1615375237
transform 1 0 2176 0 1 434
box 26 26 770 795
use cm_nmos  cm_nmos_1
timestamp 1616067151
transform 1 0 2272 0 1 6080
box -70 0 1070 4100
use en_nmos  en_nmos_0
timestamp 1616065709
transform 1 0 2272 0 1 2380
box -70 0 1070 3500
use cm_pmos  cm_pmos_0
timestamp 1616078161
transform 1 0 2272 0 1 10410
box -136 -20 1136 4100
use sky130_fd_pr__pnp_05v5_W3p40L3p40  sky130_fd_pr__pnp_05v5_W3p40L3p40_1
timestamp 1615375237
transform 1 0 2974 0 1 1250
box 26 26 770 795
use sky130_fd_pr__pnp_05v5_W3p40L3p40  sky130_fd_pr__pnp_05v5_W3p40L3p40_3
timestamp 1615375237
transform 1 0 2974 0 1 434
box 26 26 770 795
use sky130_fd_pr__pnp_05v5_W3p40L3p40  sky130_fd_pr__pnp_05v5_W3p40L3p40_6
timestamp 1615375237
transform 1 0 3772 0 1 1250
box 26 26 770 795
use sky130_fd_pr__pnp_05v5_W3p40L3p40  sky130_fd_pr__pnp_05v5_W3p40L3p40_5
timestamp 1615375237
transform 1 0 3772 0 1 434
box 26 26 770 795
use en_nmos  en_nmos_1
timestamp 1616065709
transform 1 0 3798 0 1 2380
box -70 0 1070 3500
use cm_nmos  cm_nmos_0
timestamp 1616067151
transform 1 0 3798 0 1 6080
box -70 0 1070 4100
use cm_pmos  cm_pmos_1
timestamp 1616078161
transform 1 0 3798 0 1 10410
box -136 -20 1136 4100
use sky130_fd_pr__pnp_05v5_W3p40L3p40  sky130_fd_pr__pnp_05v5_W3p40L3p40_7
timestamp 1615375237
transform 1 0 4570 0 1 1250
box 26 26 770 795
use sky130_fd_pr__pnp_05v5_W3p40L3p40  sky130_fd_pr__pnp_05v5_W3p40L3p40_4
timestamp 1615375237
transform 1 0 4570 0 1 434
box 26 26 770 795
use en_nmos  en_nmos_2
timestamp 1616065709
transform 1 0 5324 0 1 2380
box -70 0 1070 3500
use cm_pmos  cm_pmos_2
timestamp 1616078161
transform 1 0 5324 0 1 10410
box -136 -20 1136 4100
use sky130_fd_pr__pnp_05v5_W3p40L3p40  sky130_fd_pr__pnp_05v5_W3p40L3p40_8
timestamp 1615375237
transform 1 0 5368 0 1 1250
box 26 26 770 795
use sky130_fd_pr__pnp_05v5_W3p40L3p40  sky130_fd_pr__pnp_05v5_W3p40L3p40_9
timestamp 1615375237
transform 1 0 5368 0 1 434
box 26 26 770 795
<< labels >>
flabel metal1 s 6496 2226 6496 2226 0 FreeSans 400 0 0 0 A
flabel locali s 6500 5002 6500 5002 0 FreeSans 400 0 0 0 B
flabel metal1 s 4816 5982 4816 5982 0 FreeSans 400 0 0 0 C
flabel metal1 s 3768 10296 3768 10296 0 FreeSans 400 0 0 0 D
flabel metal1 s 5294 10280 5294 10280 0 FreeSans 400 0 0 0 E
flabel metal1 s 2246 2316 2246 2316 0 FreeSans 400 0 0 0 F
flabel metal1 s 3304 6000 3304 6000 0 FreeSans 400 0 0 0 G
flabel locali s 7134 11126 7134 11126 0 FreeSans 400 0 0 0 H
flabel metal1 s 7302 2132 7302 2132 0 FreeSans 400 0 0 0 J
flabel locali s 416 464 416 464 0 FreeSans 800 0 0 0 I
flabel locali s 1312 9596 1312 9596 0 FreeSans 800 0 0 0 VbiasN
flabel locali s 1628 13930 1628 13930 0 FreeSans 800 0 0 0 VbiasP
flabel locali s 404 14692 404 14692 0 FreeSans 320 0 0 0 VDD
port 0 nsew power bidirectional
flabel locali s 400 2 400 2 0 FreeSans 320 0 0 0 GND
port 1 nsew ground bidirectional
flabel locali s 7028 2336 7028 2336 0 FreeSans 320 0 0 0 Vbgp
port 2 nsew signal output
flabel locali s 6304 5360 6304 5360 0 FreeSans 320 0 0 0 en
port 3 nsew signal input
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 7636 14736
<< end >>
